/*
 *  TOPPERS/ASP Kernel
 *      Toyohashi Open Platform for Embedded Real-Time Systems/
 *      Advanced Standard Profile Kernel
 * 
 *  Copyright (C) 2015 by Ushio Laboratory
 *              Graduate School of Engineering Science, Osaka Univ., JAPAN
 *  Copyright (C) 2015,2016 by Embedded and Real-Time Systems Laboratory
 *              Graduate School of Information Science, Nagoya Univ., JAPAN
 *  Copyright (C) 2017      by Cores Co., Ltd. Japan
 * 
 *  上記著作権者は，以下の(1)～(4)の条件を満たす場合に限り，本ソフトウェ
 *  ア（本ソフトウェアを改変したものを含む．以下同じ）を使用・複製・改
 *  変・再配布（以下，利用と呼ぶ）することを無償で許諾する．
 *  (1) 本ソフトウェアをソースコードの形で利用する場合には，上記の著作
 *      権表示，この利用条件および下記の無保証規定が，そのままの形でソー
 *      スコード中に含まれていること．
 *  (2) 本ソフトウェアを，ライブラリ形式など，他のソフトウェア開発に使
 *      用できる形で再配布する場合には，再配布に伴うドキュメント（利用
 *      者マニュアルなど）に，上記の著作権表示，この利用条件および下記
 *      の無保証規定を掲載すること．
 *  (3) 本ソフトウェアを，機器に組み込むなど，他のソフトウェア開発に使
 *      用できない形で再配布する場合には，次のいずれかの条件を満たすこ
 *      と．
 *    (a) 再配布に伴うドキュメント（利用者マニュアルなど）に，上記の著
 *        作権表示，この利用条件および下記の無保証規定を掲載すること．
 *    (b) 再配布の形態を，別に定める方法によって，TOPPERSプロジェクトに
 *        報告すること．
 *  (4) 本ソフトウェアの利用により直接的または間接的に生じるいかなる損
 *      害からも，上記著作権者およびTOPPERSプロジェクトを免責すること．
 *      また，本ソフトウェアのユーザまたはエンドユーザからのいかなる理
 *      由に基づく請求からも，上記著作権者およびTOPPERSプロジェクトを
 *      免責すること．
 * 
 *  本ソフトウェアは，無保証で提供されているものである．上記著作権者お
 *  よびTOPPERSプロジェクトは，本ソフトウェアに関して，特定の使用目的
 *  に対する適合性も含めて，いかなる保証も行わない．また，本ソフトウェ
 *  アの利用により直接的または間接的に生じたいかなる損害に関しても，そ
 *  の責任を負わない．
 * 
 *  $Id$
 */

/*
 *		シリアルインタフェースドライバのターゲット依存部（GR-SAKURA用）
 *		のコンポーネント記述
 */

/*
 *  GR-SAKURAとRX631/RX63Nに関する定義
 */
import_C("gr_sakura.h");
import_C("device.h");

/*
 *  FIFO内蔵シリアルコミュニケーションインタフェース用 簡易SIOドライバ
 */
import("tMbedSerial.cdl");

/*
 *  シリアルインタフェースドライバのターゲット依存部の本体（シリアルイ
 *  ンタフェースドライバとSIOドライバを接続する部分）のセルタイプ
 */
celltype tSIOPortGRSakuraMain {
	/*
	 *  シリアルインタフェースドライバとの結合
	 */
	[inline] entry		sSIOPort	eSIOPort;
	[optional] call		siSIOCBR	ciSIOCBR;

	/*
	 *  SIOドライバとの結合
	 */
	call			sSIOPort	cSIOPort;
	[inline] entry	siSIOCBR	eiSIOCBR;
};

/*
 *  シリアルインタフェースドライバのターゲット依存部（複合コンポーネン
 *  ト）のセルタイプ
 */
composite tSIOPortGRSakura {
	/*
	 *  シリアルインタフェースドライバとの結合
	 */
	entry				sSIOPort	eSIOPort;
	[optional] call		siSIOCBR	ciSIOCBR;

	/*
	 *  属性の定義
	 */
	attr {
		int32_t tx;								/* 送信Pin */
		int32_t rx;								/* 受信Pin */
		uint32_t	baudRate = 115200;			/* ボーレートの設定値 */
	};

	/*
	 *  SIOドライバ
	 */
	cell tMbedSerial MbedSerial {
		tx          = composite.tx;
		rx          = composite.rx;
		baudRate    = composite.baudRate;
		ciSIOCBR    = SIOPortMain.eiSIOCBR;
	};

	/*
	 *  シリアルインタフェースドライバのターゲット依存部の本体
	 */
	cell tSIOPortGRSakuraMain SIOPortMain {
		ciSIOCBR            => composite.ciSIOCBR;
		cSIOPort            = MbedSerial.eSIOPort;
	};
	composite.eSIOPort => SIOPortMain.eSIOPort;
};

/*
 *  シリアルインタフェースドライバのターゲット依存部のプロトタイプ
 *
 *  サンプルプログラムが使うポートが，SIOPortTarget1に固定されているた
 *  め，ポート1とポート3を入れ換えている．具体的には，SIOPortTarget1は
 *  MbedSerialのチャネル2（チャネル番号は0から始まるので，ポート3のこと）に，
 *  SIOPortTarget3はMbedSerialのチャネル0につながっている．
 */
[prototype]
cell tSIOPortGRSakura SIOPortTarget1 {
	/* 属性の設定 */
	tx = C_EXP("P20");		/* PIN_IO1 */
	rx = C_EXP("P21");		/* PIN_IO0 */
};

[prototype]
cell tSIOPortGRSakura SIOPortTarget2 {
	/* 属性の設定 */
	tx = C_EXP("P32");		/* PIN_IO6 */
	rx = C_EXP("P33");		/* PIN_IO7 */
};

[prototype]
cell tSIOPortGRSakura SIOPortTarget3 {
	/* 属性の設定 */
	tx = C_EXP("P50");		/* PIN_IO24 */
	rx = C_EXP("P52");		/* PIN_IO26 */
};

[prototype]
cell tSIOPortGRSakura SIOPortTarget4 {
	/* 属性の設定 */
	tx = C_EXP("P23");		/* PIN_IO3 */
	rx = C_EXP("P25");		/* PIN_IO5 */
};

[prototype]
cell tSIOPortGRSakura SIOPortTarget5 {
	/* 属性の設定 */
	tx = C_EXP("PC3");		/* PIN_IO9 */
	rx = C_EXP("PC2");		/* PIN_IO8 */
};

[prototype]
cell tSIOPortGRSakura SIOPortTarget6 {
	/* 属性の設定 */
	tx = C_EXP("PC7");		/* PIN_IO12 */
	rx = C_EXP("PC6");		/* PIN_IO11 */
};

[prototype]
cell tSIOPortGRSakura SIOPortTarget7 {
	/* 属性の設定 */
	tx = C_EXP("P26");		/* PIN_IO58 */
	rx = C_EXP("P30");		/* PIN_IO60 */
};

[prototype]
cell tSIOPortGRSakura SIOPortTarget8 {
	/* 属性の設定 */
	tx = NULL;
	rx = NULL;
};
